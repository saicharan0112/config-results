module tempsenseInst_error (CLK_REF,
    DONE,
    RESET_COUNTERn,
    en,
    lc_out,
    out,
    outb,
    \r_VIN(0) ,
    \r_VIN(1) ,
    \r_VIN(2) ,
    DOUT,
    SEL_CONV_TIME);
 input CLK_REF;
 output DONE;
 input RESET_COUNTERn;
 input en;
 output lc_out;
 output out;
 output outb;
 input \r_VIN(0) ;
 input \r_VIN(1) ;
 input \r_VIN(2) ;
 output [23:0] DOUT;
 input [3:0] SEL_CONV_TIME;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _067_;
 wire _068_;
 wire \temp_analog_0.n1 ;
 wire \temp_analog_0.n2 ;
 wire \temp_analog_0.n3 ;
 wire \temp_analog_0.n4 ;
 wire \temp_analog_0.n5 ;
 wire \temp_analog_0.n6 ;
 wire \temp_analog_0.n7 ;
 wire r_VIN;
 wire \temp_analog_0.nx2 ;
 wire \temp_analog_1.VIN ;
 wire \temp_analog_1.async_counter_0.WAKE ;
 wire \temp_analog_1.async_counter_0.WAKE_pre ;
 wire \temp_analog_1.async_counter_0.clk_ref_in ;
 wire \temp_analog_1.async_counter_0.clk_sens_in ;
 wire \temp_analog_1.async_counter_0.div_r[0] ;
 wire \temp_analog_1.async_counter_0.div_r[10] ;
 wire \temp_analog_1.async_counter_0.div_r[11] ;
 wire \temp_analog_1.async_counter_0.div_r[12] ;
 wire \temp_analog_1.async_counter_0.div_r[13] ;
 wire \temp_analog_1.async_counter_0.div_r[14] ;
 wire \temp_analog_1.async_counter_0.div_r[15] ;
 wire \temp_analog_1.async_counter_0.div_r[16] ;
 wire \temp_analog_1.async_counter_0.div_r[17] ;
 wire \temp_analog_1.async_counter_0.div_r[18] ;
 wire \temp_analog_1.async_counter_0.div_r[19] ;
 wire \temp_analog_1.async_counter_0.div_r[1] ;
 wire \temp_analog_1.async_counter_0.div_r[20] ;
 wire \temp_analog_1.async_counter_0.div_r[2] ;
 wire \temp_analog_1.async_counter_0.div_r[3] ;
 wire \temp_analog_1.async_counter_0.div_r[4] ;
 wire \temp_analog_1.async_counter_0.div_r[5] ;
 wire \temp_analog_1.async_counter_0.div_r[6] ;
 wire \temp_analog_1.async_counter_0.div_r[7] ;
 wire \temp_analog_1.async_counter_0.div_r[8] ;
 wire \temp_analog_1.async_counter_0.div_r[9] ;
 wire \temp_analog_1.async_counter_0.div_s[0] ;
 wire \temp_analog_1.async_counter_0.div_s[10] ;
 wire \temp_analog_1.async_counter_0.div_s[11] ;
 wire \temp_analog_1.async_counter_0.div_s[12] ;
 wire \temp_analog_1.async_counter_0.div_s[13] ;
 wire \temp_analog_1.async_counter_0.div_s[14] ;
 wire \temp_analog_1.async_counter_0.div_s[15] ;
 wire \temp_analog_1.async_counter_0.div_s[16] ;
 wire \temp_analog_1.async_counter_0.div_s[17] ;
 wire \temp_analog_1.async_counter_0.div_s[18] ;
 wire \temp_analog_1.async_counter_0.div_s[19] ;
 wire \temp_analog_1.async_counter_0.div_s[1] ;
 wire \temp_analog_1.async_counter_0.div_s[20] ;
 wire \temp_analog_1.async_counter_0.div_s[21] ;
 wire \temp_analog_1.async_counter_0.div_s[22] ;
 wire \temp_analog_1.async_counter_0.div_s[23] ;
 wire \temp_analog_1.async_counter_0.div_s[2] ;
 wire \temp_analog_1.async_counter_0.div_s[3] ;
 wire \temp_analog_1.async_counter_0.div_s[4] ;
 wire \temp_analog_1.async_counter_0.div_s[5] ;
 wire \temp_analog_1.async_counter_0.div_s[6] ;
 wire \temp_analog_1.async_counter_0.div_s[7] ;
 wire \temp_analog_1.async_counter_0.div_s[8] ;
 wire \temp_analog_1.async_counter_0.div_s[9] ;

 sky130_fd_sc_hd__inv_1 _069_ (.A(\temp_analog_1.async_counter_0.div_r[5] ),
    .Y(_068_));
 sky130_fd_sc_hd__inv_1 _070_ (.A(\temp_analog_1.async_counter_0.div_r[19] ),
    .Y(_036_));
 sky130_fd_sc_hd__inv_1 _071_ (.A(\temp_analog_1.async_counter_0.div_r[18] ),
    .Y(_037_));
 sky130_fd_sc_hd__inv_1 _072_ (.A(\temp_analog_1.async_counter_0.div_r[17] ),
    .Y(_038_));
 sky130_fd_sc_hd__inv_1 _073_ (.A(\temp_analog_1.async_counter_0.div_r[16] ),
    .Y(_039_));
 sky130_fd_sc_hd__inv_1 _074_ (.A(\temp_analog_1.async_counter_0.div_r[15] ),
    .Y(_040_));
 sky130_fd_sc_hd__inv_1 _075_ (.A(\temp_analog_1.async_counter_0.div_r[14] ),
    .Y(_041_));
 sky130_fd_sc_hd__inv_1 _076_ (.A(\temp_analog_1.async_counter_0.div_r[13] ),
    .Y(_042_));
 sky130_fd_sc_hd__inv_1 _077_ (.A(\temp_analog_1.async_counter_0.div_r[12] ),
    .Y(_043_));
 sky130_fd_sc_hd__inv_1 _078_ (.A(\temp_analog_1.async_counter_0.div_r[11] ),
    .Y(_044_));
 sky130_fd_sc_hd__inv_1 _079_ (.A(\temp_analog_1.async_counter_0.div_r[10] ),
    .Y(_031_));
 sky130_fd_sc_hd__inv_1 _080_ (.A(\temp_analog_1.async_counter_0.div_r[9] ),
    .Y(_032_));
 sky130_fd_sc_hd__inv_1 _081_ (.A(\temp_analog_1.async_counter_0.div_r[8] ),
    .Y(_033_));
 sky130_fd_sc_hd__inv_1 _082_ (.A(\temp_analog_1.async_counter_0.div_r[7] ),
    .Y(_034_));
 sky130_fd_sc_hd__inv_1 _083_ (.A(\temp_analog_1.async_counter_0.div_r[6] ),
    .Y(_035_));
 sky130_fd_sc_hd__inv_1 _084_ (.A(SEL_CONV_TIME[3]),
    .Y(_045_));
 sky130_fd_sc_hd__decap_4 PHY_12 ();
 sky130_fd_sc_hd__decap_4 PHY_11 ();
 sky130_fd_sc_hd__nor3_1 _087_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(\temp_analog_1.async_counter_0.div_r[17] ),
    .Y(_048_));
 sky130_fd_sc_hd__or2b_1 _088_ (.A(SEL_CONV_TIME[0]),
    .B_N(SEL_CONV_TIME[1]),
    .X(_049_));
 sky130_fd_sc_hd__nand2_1 _089_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .Y(_050_));
 sky130_fd_sc_hd__or3b_2 _090_ (.A(SEL_CONV_TIME[1]),
    .B(\temp_analog_1.async_counter_0.div_r[18] ),
    .C_N(SEL_CONV_TIME[0]),
    .X(_051_));
 sky130_fd_sc_hd__o221ai_1 _091_ (.A1(\temp_analog_1.async_counter_0.div_r[19] ),
    .A2(_049_),
    .B1(_050_),
    .B2(\temp_analog_1.async_counter_0.div_r[20] ),
    .C1(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__mux4_1 _092_ (.A0(\temp_analog_1.async_counter_0.div_r[9] ),
    .A1(\temp_analog_1.async_counter_0.div_r[10] ),
    .A2(\temp_analog_1.async_counter_0.div_r[11] ),
    .A3(\temp_analog_1.async_counter_0.div_r[12] ),
    .S0(SEL_CONV_TIME[0]),
    .S1(SEL_CONV_TIME[1]),
    .X(_053_));
 sky130_fd_sc_hd__nand2_1 _093_ (.A(_045_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__o311a_1 _094_ (.A1(_045_),
    .A2(_048_),
    .A3(_052_),
    .B1(_054_),
    .C1(SEL_CONV_TIME[2]),
    .X(_055_));
 sky130_fd_sc_hd__decap_4 PHY_10 ();
 sky130_fd_sc_hd__nand3b_1 _096_ (.A_N(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(_041_),
    .Y(_057_));
 sky130_fd_sc_hd__or3_1 _097_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(\temp_analog_1.async_counter_0.div_r[13] ),
    .X(_058_));
 sky130_fd_sc_hd__nand3b_1 _098_ (.A_N(\temp_analog_1.async_counter_0.div_r[16] ),
    .B(SEL_CONV_TIME[0]),
    .C(SEL_CONV_TIME[1]),
    .Y(_059_));
 sky130_fd_sc_hd__o2111a_2 _099_ (.A1(\temp_analog_1.async_counter_0.div_r[15] ),
    .A2(_049_),
    .B1(_058_),
    .C1(_059_),
    .D1(SEL_CONV_TIME[3]),
    .X(_060_));
 sky130_fd_sc_hd__mux4_2 _100_ (.A0(\temp_analog_1.async_counter_0.div_r[5] ),
    .A1(\temp_analog_1.async_counter_0.div_r[7] ),
    .A2(\temp_analog_1.async_counter_0.div_r[6] ),
    .A3(\temp_analog_1.async_counter_0.div_r[8] ),
    .S0(SEL_CONV_TIME[1]),
    .S1(SEL_CONV_TIME[0]),
    .X(_061_));
 sky130_fd_sc_hd__a221oi_4 _101_ (.A1(_057_),
    .A2(_060_),
    .B1(_061_),
    .B2(_045_),
    .C1(SEL_CONV_TIME[2]),
    .Y(_062_));
 sky130_fd_sc_hd__o211a_1 _102_ (.A1(_055_),
    .A2(_062_),
    .B1(\temp_analog_1.async_counter_0.WAKE ),
    .C1(CLK_REF),
    .X(\temp_analog_1.async_counter_0.clk_ref_in ));
 sky130_fd_sc_hd__o211a_1 _103_ (.A1(_055_),
    .A2(_062_),
    .B1(\temp_analog_1.async_counter_0.WAKE_pre ),
    .C1(lc_out),
    .X(\temp_analog_1.async_counter_0.clk_sens_in ));
 sky130_fd_sc_hd__inv_1 _104_ (.A(\temp_analog_1.async_counter_0.div_s[0] ),
    .Y(_005_));
 sky130_fd_sc_hd__decap_4 PHY_9 ();
 sky130_fd_sc_hd__decap_4 PHY_8 ();
 sky130_fd_sc_hd__nor3_2 _107_ (.A(_005_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[0]));
 sky130_fd_sc_hd__inv_1 _108_ (.A(\temp_analog_1.async_counter_0.div_s[1] ),
    .Y(_016_));
 sky130_fd_sc_hd__nor3_2 _109_ (.A(_016_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[1]));
 sky130_fd_sc_hd__inv_1 _110_ (.A(\temp_analog_1.async_counter_0.div_s[2] ),
    .Y(_021_));
 sky130_fd_sc_hd__nor3_2 _111_ (.A(_021_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[2]));
 sky130_fd_sc_hd__inv_1 _112_ (.A(\temp_analog_1.async_counter_0.div_s[3] ),
    .Y(_022_));
 sky130_fd_sc_hd__nor3_1 _113_ (.A(_022_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[3]));
 sky130_fd_sc_hd__inv_1 _114_ (.A(\temp_analog_1.async_counter_0.div_s[4] ),
    .Y(_023_));
 sky130_fd_sc_hd__nor3_2 _115_ (.A(_023_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[4]));
 sky130_fd_sc_hd__inv_1 _116_ (.A(\temp_analog_1.async_counter_0.div_s[5] ),
    .Y(_024_));
 sky130_fd_sc_hd__nor3_1 _117_ (.A(_024_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[5]));
 sky130_fd_sc_hd__inv_1 _118_ (.A(\temp_analog_1.async_counter_0.div_s[6] ),
    .Y(_025_));
 sky130_fd_sc_hd__nor3_1 _119_ (.A(_025_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[6]));
 sky130_fd_sc_hd__inv_1 _120_ (.A(\temp_analog_1.async_counter_0.div_s[7] ),
    .Y(_026_));
 sky130_fd_sc_hd__nor3_1 _121_ (.A(_026_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[7]));
 sky130_fd_sc_hd__inv_1 _122_ (.A(\temp_analog_1.async_counter_0.div_s[8] ),
    .Y(_027_));
 sky130_fd_sc_hd__nor3_1 _123_ (.A(_027_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[8]));
 sky130_fd_sc_hd__inv_1 _124_ (.A(\temp_analog_1.async_counter_0.div_s[9] ),
    .Y(_028_));
 sky130_fd_sc_hd__decap_4 PHY_7 ();
 sky130_fd_sc_hd__decap_4 PHY_6 ();
 sky130_fd_sc_hd__nor3_1 _127_ (.A(_028_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[9]));
 sky130_fd_sc_hd__inv_1 _128_ (.A(\temp_analog_1.async_counter_0.div_s[10] ),
    .Y(_006_));
 sky130_fd_sc_hd__nor3_1 _129_ (.A(_006_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[10]));
 sky130_fd_sc_hd__inv_1 _130_ (.A(\temp_analog_1.async_counter_0.div_s[11] ),
    .Y(_007_));
 sky130_fd_sc_hd__nor3_1 _131_ (.A(_007_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[11]));
 sky130_fd_sc_hd__inv_1 _132_ (.A(\temp_analog_1.async_counter_0.div_s[12] ),
    .Y(_008_));
 sky130_fd_sc_hd__nor3_1 _133_ (.A(_008_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[12]));
 sky130_fd_sc_hd__inv_1 _134_ (.A(\temp_analog_1.async_counter_0.div_s[13] ),
    .Y(_009_));
 sky130_fd_sc_hd__nor3_1 _135_ (.A(_009_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[13]));
 sky130_fd_sc_hd__inv_1 _136_ (.A(\temp_analog_1.async_counter_0.div_s[14] ),
    .Y(_010_));
 sky130_fd_sc_hd__nor3_1 _137_ (.A(_010_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[14]));
 sky130_fd_sc_hd__inv_1 _138_ (.A(\temp_analog_1.async_counter_0.div_s[15] ),
    .Y(_011_));
 sky130_fd_sc_hd__nor3_1 _139_ (.A(_011_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[15]));
 sky130_fd_sc_hd__inv_1 _140_ (.A(\temp_analog_1.async_counter_0.div_s[16] ),
    .Y(_012_));
 sky130_fd_sc_hd__nor3_1 _141_ (.A(_012_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[16]));
 sky130_fd_sc_hd__inv_1 _142_ (.A(\temp_analog_1.async_counter_0.div_s[17] ),
    .Y(_013_));
 sky130_fd_sc_hd__nor3_1 _143_ (.A(_013_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[17]));
 sky130_fd_sc_hd__inv_1 _144_ (.A(\temp_analog_1.async_counter_0.div_s[18] ),
    .Y(_014_));
 sky130_fd_sc_hd__nor3_1 _145_ (.A(_014_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[18]));
 sky130_fd_sc_hd__inv_1 _146_ (.A(\temp_analog_1.async_counter_0.div_s[19] ),
    .Y(_015_));
 sky130_fd_sc_hd__nor3_1 _147_ (.A(_015_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[19]));
 sky130_fd_sc_hd__inv_1 _148_ (.A(\temp_analog_1.async_counter_0.div_s[20] ),
    .Y(_017_));
 sky130_fd_sc_hd__nor3_1 _149_ (.A(_017_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[20]));
 sky130_fd_sc_hd__inv_1 _150_ (.A(\temp_analog_1.async_counter_0.div_s[21] ),
    .Y(_018_));
 sky130_fd_sc_hd__nor3_1 _151_ (.A(_018_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[21]));
 sky130_fd_sc_hd__inv_1 _152_ (.A(\temp_analog_1.async_counter_0.div_s[22] ),
    .Y(_019_));
 sky130_fd_sc_hd__nor3_1 _153_ (.A(_019_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[22]));
 sky130_fd_sc_hd__inv_1 _154_ (.A(\temp_analog_1.async_counter_0.div_s[23] ),
    .Y(_020_));
 sky130_fd_sc_hd__nor3_1 _155_ (.A(_020_),
    .B(_055_),
    .C(_062_),
    .Y(DOUT[23]));
 sky130_fd_sc_hd__nor2_1 _156_ (.A(_055_),
    .B(_062_),
    .Y(DONE));
 sky130_fd_sc_hd__inv_1 _157_ (.A(\temp_analog_1.async_counter_0.div_r[20] ),
    .Y(_030_));
 sky130_fd_sc_hd__inv_1 _158_ (.A(\temp_analog_1.async_counter_0.div_r[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_1 _159_ (.A(\temp_analog_1.async_counter_0.div_r[1] ),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _160_ (.A(\temp_analog_1.async_counter_0.div_r[2] ),
    .Y(_002_));
 sky130_fd_sc_hd__inv_1 _161_ (.A(\temp_analog_1.async_counter_0.div_r[3] ),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _162_ (.A(\temp_analog_1.async_counter_0.div_r[4] ),
    .Y(_004_));
 sky130_fd_sc_hd__or2_2 _163_ (.A(\temp_analog_1.async_counter_0.WAKE ),
    .B(\temp_analog_1.async_counter_0.WAKE_pre ),
    .X(_029_));
 sky130_fd_sc_hd__dfrtp_1 _164_ (.D(_029_),
    .Q(\temp_analog_1.async_counter_0.WAKE ),
    .RESET_B(RESET_COUNTERn),
    .CLK(CLK_REF));
 sky130_fd_sc_hd__dfrtp_1 _165_ (.D(_067_),
    .Q(\temp_analog_1.async_counter_0.WAKE_pre ),
    .RESET_B(RESET_COUNTERn),
    .CLK(CLK_REF));
 sky130_fd_sc_hd__dfrtn_1 _166_ (.D(_030_),
    .Q(\temp_analog_1.async_counter_0.div_r[20] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[19] ));
 sky130_fd_sc_hd__dfrtn_1 _167_ (.D(_036_),
    .Q(\temp_analog_1.async_counter_0.div_r[19] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[18] ));
 sky130_fd_sc_hd__dfrtn_1 _168_ (.D(_037_),
    .Q(\temp_analog_1.async_counter_0.div_r[18] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[17] ));
 sky130_fd_sc_hd__dfrtn_1 _169_ (.D(_038_),
    .Q(\temp_analog_1.async_counter_0.div_r[17] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[16] ));
 sky130_fd_sc_hd__dfrtn_1 _170_ (.D(_039_),
    .Q(\temp_analog_1.async_counter_0.div_r[16] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[15] ));
 sky130_fd_sc_hd__dfrtn_1 _171_ (.D(_040_),
    .Q(\temp_analog_1.async_counter_0.div_r[15] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[14] ));
 sky130_fd_sc_hd__dfrtn_1 _172_ (.D(_041_),
    .Q(\temp_analog_1.async_counter_0.div_r[14] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[13] ));
 sky130_fd_sc_hd__dfrtn_1 _173_ (.D(_042_),
    .Q(\temp_analog_1.async_counter_0.div_r[13] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[12] ));
 sky130_fd_sc_hd__dfrtn_1 _174_ (.D(_043_),
    .Q(\temp_analog_1.async_counter_0.div_r[12] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[11] ));
 sky130_fd_sc_hd__dfrtn_1 _175_ (.D(_044_),
    .Q(\temp_analog_1.async_counter_0.div_r[11] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[10] ));
 sky130_fd_sc_hd__dfrtn_1 _176_ (.D(_031_),
    .Q(\temp_analog_1.async_counter_0.div_r[10] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[9] ));
 sky130_fd_sc_hd__dfrtn_1 _177_ (.D(_032_),
    .Q(\temp_analog_1.async_counter_0.div_r[9] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[8] ));
 sky130_fd_sc_hd__dfrtn_1 _178_ (.D(_033_),
    .Q(\temp_analog_1.async_counter_0.div_r[8] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[7] ));
 sky130_fd_sc_hd__dfrtn_1 _179_ (.D(_034_),
    .Q(\temp_analog_1.async_counter_0.div_r[7] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[6] ));
 sky130_fd_sc_hd__dfrtn_1 _180_ (.D(_035_),
    .Q(\temp_analog_1.async_counter_0.div_r[6] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[5] ));
 sky130_fd_sc_hd__dfrtn_1 _181_ (.D(_068_),
    .Q(\temp_analog_1.async_counter_0.div_r[5] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[4] ));
 sky130_fd_sc_hd__dfrtn_1 _182_ (.D(_004_),
    .Q(\temp_analog_1.async_counter_0.div_r[4] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[3] ));
 sky130_fd_sc_hd__dfrtn_1 _183_ (.D(_003_),
    .Q(\temp_analog_1.async_counter_0.div_r[3] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[2] ));
 sky130_fd_sc_hd__dfrtn_1 _184_ (.D(_002_),
    .Q(\temp_analog_1.async_counter_0.div_r[2] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[1] ));
 sky130_fd_sc_hd__dfrtn_1 _185_ (.D(_001_),
    .Q(\temp_analog_1.async_counter_0.div_r[1] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_r[0] ));
 sky130_fd_sc_hd__dfrtn_1 _186_ (.D(_020_),
    .Q(\temp_analog_1.async_counter_0.div_s[23] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[22] ));
 sky130_fd_sc_hd__dfrtn_1 _187_ (.D(_019_),
    .Q(\temp_analog_1.async_counter_0.div_s[22] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[21] ));
 sky130_fd_sc_hd__dfrtn_1 _188_ (.D(_018_),
    .Q(\temp_analog_1.async_counter_0.div_s[21] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[20] ));
 sky130_fd_sc_hd__dfrtn_1 _189_ (.D(_017_),
    .Q(\temp_analog_1.async_counter_0.div_s[20] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[19] ));
 sky130_fd_sc_hd__dfrtn_1 _190_ (.D(_015_),
    .Q(\temp_analog_1.async_counter_0.div_s[19] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[18] ));
 sky130_fd_sc_hd__dfrtn_1 _191_ (.D(_014_),
    .Q(\temp_analog_1.async_counter_0.div_s[18] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[17] ));
 sky130_fd_sc_hd__dfrtn_1 _192_ (.D(_013_),
    .Q(\temp_analog_1.async_counter_0.div_s[17] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[16] ));
 sky130_fd_sc_hd__dfrtn_1 _193_ (.D(_012_),
    .Q(\temp_analog_1.async_counter_0.div_s[16] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[15] ));
 sky130_fd_sc_hd__dfrtn_1 _194_ (.D(_011_),
    .Q(\temp_analog_1.async_counter_0.div_s[15] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[14] ));
 sky130_fd_sc_hd__dfrtn_1 _195_ (.D(_010_),
    .Q(\temp_analog_1.async_counter_0.div_s[14] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[13] ));
 sky130_fd_sc_hd__dfrtn_1 _196_ (.D(_009_),
    .Q(\temp_analog_1.async_counter_0.div_s[13] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[12] ));
 sky130_fd_sc_hd__dfrtn_1 _197_ (.D(_008_),
    .Q(\temp_analog_1.async_counter_0.div_s[12] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[11] ));
 sky130_fd_sc_hd__dfrtn_1 _198_ (.D(_007_),
    .Q(\temp_analog_1.async_counter_0.div_s[11] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[10] ));
 sky130_fd_sc_hd__dfrtn_1 _199_ (.D(_006_),
    .Q(\temp_analog_1.async_counter_0.div_s[10] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[9] ));
 sky130_fd_sc_hd__dfrtn_1 _200_ (.D(_028_),
    .Q(\temp_analog_1.async_counter_0.div_s[9] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[8] ));
 sky130_fd_sc_hd__dfrtn_1 _201_ (.D(_027_),
    .Q(\temp_analog_1.async_counter_0.div_s[8] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[7] ));
 sky130_fd_sc_hd__dfrtn_1 _202_ (.D(_026_),
    .Q(\temp_analog_1.async_counter_0.div_s[7] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[6] ));
 sky130_fd_sc_hd__dfrtn_1 _203_ (.D(_025_),
    .Q(\temp_analog_1.async_counter_0.div_s[6] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[5] ));
 sky130_fd_sc_hd__dfrtn_1 _204_ (.D(_024_),
    .Q(\temp_analog_1.async_counter_0.div_s[5] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[4] ));
 sky130_fd_sc_hd__dfrtn_1 _205_ (.D(_023_),
    .Q(\temp_analog_1.async_counter_0.div_s[4] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[3] ));
 sky130_fd_sc_hd__dfrtn_1 _206_ (.D(_022_),
    .Q(\temp_analog_1.async_counter_0.div_s[3] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[2] ));
 sky130_fd_sc_hd__dfrtn_1 _207_ (.D(_021_),
    .Q(\temp_analog_1.async_counter_0.div_s[2] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[1] ));
 sky130_fd_sc_hd__dfrtn_1 _208_ (.D(_016_),
    .Q(\temp_analog_1.async_counter_0.div_s[1] ),
    .RESET_B(RESET_COUNTERn),
    .CLK_N(\temp_analog_1.async_counter_0.div_s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _209_ (.D(_000_),
    .Q(\temp_analog_1.async_counter_0.div_r[0] ),
    .RESET_B(RESET_COUNTERn),
    .CLK(\temp_analog_1.async_counter_0.clk_ref_in ));
 sky130_fd_sc_hd__dfrtp_1 _210_ (.D(_005_),
    .Q(\temp_analog_1.async_counter_0.div_s[0] ),
    .RESET_B(RESET_COUNTERn),
    .CLK(\temp_analog_1.async_counter_0.clk_sens_in ));
 sky130_fd_sc_hd__conb_1 _211_ (.HI(_067_));
 sky130_fd_sc_hd__decap_4 PHY_5 ();
 sky130_fd_sc_hd__decap_4 PHY_4 ();
 sky130_fd_sc_hd__decap_4 PHY_3 ();
 sky130_fd_sc_hd__decap_4 PHY_2 ();
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_0  (.A(\temp_analog_0.n1 ),
    .Y(\temp_analog_0.n2 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_1  (.A(\temp_analog_0.n2 ),
    .Y(\temp_analog_0.n3 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_2  (.A(\temp_analog_0.n3 ),
    .Y(\temp_analog_0.n4 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_3  (.A(\temp_analog_0.n4 ),
    .Y(\temp_analog_0.n5 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_4  (.A(\temp_analog_0.n5 ),
    .Y(\temp_analog_0.n6 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_5  (.A(\temp_analog_0.n6 ),
    .Y(\temp_analog_0.n7 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m1  (.A(\temp_analog_0.n7 ),
    .Y(out));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m2  (.A(\temp_analog_0.n7 ),
    .Y(\temp_analog_0.nx2 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m3  (.A(\temp_analog_0.nx2 ),
    .Y(outb));
 sky130_fd_sc_hd__nand2_1 \temp_analog_0.a_nand_0  (.A(en),
    .B(\temp_analog_0.n7 ),
    .Y(\temp_analog_0.n1 ));
 sky130_fd_sc_hd__decap_4 PHY_1 ();
 HEADER \temp_analog_1.a_header_0  (.VIN(r_VIN));
 HEADER \temp_analog_1.a_header_1  (.VIN(r_VIN));
 HEADER \temp_analog_1.a_header_2  (.VIN(r_VIN));
 HEADER \temp_analog_1.a_header_3  (.VIN(r_VIN));
 HEADER \temp_analog_1.a_header_4  (.VIN(r_VIN));
 SLC \temp_analog_1.a_lc_0  (.IN(out),
    .INB(outb),
    .VOUT(lc_out));
 sky130_fd_sc_hd__decap_4 PHY_0 ();
 sky130_fd_sc_hd__decap_4 PHY_13 ();
 sky130_fd_sc_hd__decap_4 PHY_14 ();
 sky130_fd_sc_hd__decap_4 PHY_15 ();
 sky130_fd_sc_hd__decap_4 PHY_16 ();
 sky130_fd_sc_hd__decap_4 PHY_17 ();
 sky130_fd_sc_hd__decap_4 PHY_18 ();
 sky130_fd_sc_hd__decap_4 PHY_19 ();
 sky130_fd_sc_hd__decap_4 PHY_20 ();
 sky130_fd_sc_hd__decap_4 PHY_21 ();
 sky130_fd_sc_hd__decap_4 PHY_22 ();
 sky130_fd_sc_hd__decap_4 PHY_23 ();
 sky130_fd_sc_hd__decap_4 PHY_24 ();
 sky130_fd_sc_hd__decap_4 PHY_25 ();
 sky130_fd_sc_hd__decap_4 PHY_26 ();
 sky130_fd_sc_hd__decap_4 PHY_27 ();
 sky130_fd_sc_hd__decap_4 PHY_28 ();
 sky130_fd_sc_hd__decap_4 PHY_29 ();
 sky130_fd_sc_hd__decap_4 PHY_30 ();
 sky130_fd_sc_hd__decap_4 PHY_31 ();
 sky130_fd_sc_hd__decap_4 PHY_32 ();
 sky130_fd_sc_hd__decap_4 PHY_33 ();
 sky130_fd_sc_hd__decap_4 PHY_34 ();
 sky130_fd_sc_hd__decap_4 PHY_35 ();
 sky130_fd_sc_hd__decap_4 PHY_36 ();
 sky130_fd_sc_hd__decap_4 PHY_37 ();
 sky130_fd_sc_hd__decap_4 PHY_38 ();
 sky130_fd_sc_hd__decap_4 PHY_39 ();
 sky130_fd_sc_hd__decap_4 PHY_40 ();
 sky130_fd_sc_hd__decap_4 PHY_41 ();
 sky130_fd_sc_hd__decap_4 PHY_42 ();
 sky130_fd_sc_hd__decap_4 PHY_43 ();
 sky130_fd_sc_hd__decap_4 PHY_44 ();
 sky130_fd_sc_hd__decap_4 PHY_45 ();
 sky130_fd_sc_hd__decap_4 PHY_46 ();
 sky130_fd_sc_hd__decap_4 PHY_47 ();
 sky130_fd_sc_hd__decap_4 PHY_48 ();
 sky130_fd_sc_hd__decap_4 PHY_49 ();
 sky130_fd_sc_hd__decap_4 PHY_50 ();
 sky130_fd_sc_hd__decap_4 PHY_51 ();
 sky130_fd_sc_hd__decap_4 PHY_52 ();
 sky130_fd_sc_hd__decap_4 PHY_53 ();
 sky130_fd_sc_hd__decap_4 PHY_54 ();
 sky130_fd_sc_hd__decap_4 PHY_55 ();
 sky130_fd_sc_hd__decap_4 PHY_56 ();
 sky130_fd_sc_hd__decap_4 PHY_57 ();
 sky130_fd_sc_hd__decap_4 PHY_58 ();
 sky130_fd_sc_hd__decap_4 PHY_59 ();
 sky130_fd_sc_hd__decap_4 PHY_60 ();
 sky130_fd_sc_hd__decap_4 PHY_61 ();
 sky130_fd_sc_hd__decap_4 PHY_62 ();
 sky130_fd_sc_hd__decap_4 PHY_63 ();
 sky130_fd_sc_hd__decap_4 PHY_64 ();
 sky130_fd_sc_hd__decap_4 PHY_65 ();
 sky130_fd_sc_hd__decap_4 PHY_66 ();
 sky130_fd_sc_hd__decap_4 PHY_67 ();
 sky130_fd_sc_hd__decap_4 PHY_68 ();
 sky130_fd_sc_hd__decap_4 PHY_69 ();
 sky130_fd_sc_hd__decap_4 PHY_70 ();
 sky130_fd_sc_hd__decap_4 PHY_71 ();
 sky130_fd_sc_hd__decap_4 PHY_72 ();
 sky130_fd_sc_hd__decap_4 PHY_73 ();
 sky130_fd_sc_hd__decap_4 PHY_74 ();
 sky130_fd_sc_hd__decap_4 PHY_75 ();
 sky130_fd_sc_hd__decap_4 PHY_76 ();
 sky130_fd_sc_hd__decap_4 PHY_77 ();
 sky130_fd_sc_hd__decap_4 PHY_78 ();
 sky130_fd_sc_hd__decap_4 PHY_79 ();
 sky130_fd_sc_hd__decap_4 PHY_80 ();
 sky130_fd_sc_hd__decap_4 PHY_81 ();
 sky130_fd_sc_hd__decap_4 PHY_82 ();
 sky130_fd_sc_hd__decap_4 PHY_83 ();
 sky130_fd_sc_hd__decap_4 PHY_84 ();
 sky130_fd_sc_hd__decap_4 PHY_85 ();
 sky130_fd_sc_hd__decap_4 PHY_86 ();
 sky130_fd_sc_hd__decap_4 PHY_87 ();
 sky130_fd_sc_hd__decap_4 PHY_88 ();
 sky130_fd_sc_hd__decap_4 PHY_89 ();
 sky130_fd_sc_hd__decap_4 PHY_90 ();
 sky130_fd_sc_hd__decap_4 PHY_91 ();
 sky130_fd_sc_hd__decap_4 PHY_92 ();
 sky130_fd_sc_hd__decap_4 PHY_93 ();
 sky130_fd_sc_hd__decap_4 PHY_94 ();
 sky130_fd_sc_hd__decap_4 PHY_95 ();
 sky130_fd_sc_hd__decap_4 PHY_96 ();
 sky130_fd_sc_hd__decap_4 PHY_97 ();
 sky130_fd_sc_hd__decap_4 PHY_98 ();
 sky130_fd_sc_hd__decap_4 PHY_99 ();
 sky130_fd_sc_hd__decap_4 PHY_100 ();
 sky130_fd_sc_hd__decap_4 PHY_101 ();
 sky130_fd_sc_hd__decap_4 PHY_102 ();
 sky130_fd_sc_hd__decap_4 PHY_103 ();
 sky130_fd_sc_hd__decap_4 PHY_104 ();
 sky130_fd_sc_hd__decap_4 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_253 ();
endmodule
